module CAND(
	input br,zf,
	output compand
);


assign compand=br & zf;
endmodule
