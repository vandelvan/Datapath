module MUX5(
	input [7:0] add1,
	input compand,
	output reg [7:0] pc
);

always @*
	begin
		if(compand)
		begin
			pc=add1;//iria ALUresult
		end
		else
		begin
			pc=add1;
		end
	end
endmodule
